module graytb;
reg [3:0] B;
wire [3:0] G;
graycon g1(B,G);
initial
begin
/*B[3] = 1'b0; B[2] = 1'b0; B[1] = 1'b0; B[0] = 1'b0; #5;
B[3] = 1'b0; B[2] = 1'b0; B[1] = 1'b0; B[0] = 1'b1; #5;
B[3] = 1'b0; B[2] = 1'b0; B[1] = 1'b1; B[0] = 1'b0; #5;
B[3] = 1'b0; B[2] = 1'b0; B[1] = 1'b1; B[0] = 1'b1; #5;
B[3] = 1'b0; B[2] = 1'b1; B[1] = 1'b0; B[0] = 1'b0; #5;
B[3] = 1'b0; B[2] = 1'b1; B[1] = 1'b0; B[0] = 1'b1; #5;
B[3] = 1'b0; B[2] = 1'b1; B[1] = 1'b1; B[0] = 1'b0; #5;
B[3] = 1'b0; B[2] = 1'b1; B[1] = 1'b1; B[0] = 1'b1; #5;
B[3] = 1'b1; B[2] = 1'b0; B[1] = 1'b0; B[0] = 1'b0; #5;
B[3] = 1'b1; B[2] = 1'b0; B[1] = 1'b0; B[0] = 1'b1; #5;
B[3] = 1'b1; B[2] = 1'b0; B[1] = 1'b1; B[0] = 1'b0; #5;
B[3] = 1'b1; B[2] = 1'b0; B[1] = 1'b1; B[0] = 1'b1; #5;
B[3] = 1'b1; B[2] = 1'b1; B[1] = 1'b0; B[0] = 1'b0; #5;
B[3] = 1'b1; B[2] = 1'b1; B[1] = 1'b0; B[0] = 1'b1; #5;
B[3] = 1'b1; B[2] = 1'b1; B[1] = 1'b1; B[0] = 1'b0; #5;
B[3] = 1'b1; B[2] = 1'b1; B[1] = 1'b1; B[0] = 1'b1; #5;*/
B=4'b0000; #5
B=4'b0001; #5
B=4'b0011; #5
B=4'b0111; #5;

end
endmodule;
